`timescale 1ns/1ns
`include "dec4_16.v"

module dec4_16_tb;

reg a,b,c,d;
output [15:0] o;

dec4_16 uut(a,b,c,d,o);

initial begin
    
    $dumpfile("dec4_16_tb.vcd");
    $dumpvars(0 , dec4_16_tb);

    a = 0; b = 0; c = 0; d = 0; #10;
    a = 0; b = 0; c = 0; d = 1; #10;
    a = 0; b = 0; c = 1; d = 0; #10;
    a = 0; b = 0; c = 1; d = 1; #10;
    a = 0; b = 1; c = 0; d = 0; #10;
    a = 0; b = 1; c = 0; d = 1; #10;
    a = 0; b = 1; c = 1; d = 0; #10;
    a = 0; b = 1; c = 1; d = 1; #10;
    a = 1; b = 0; c = 0; d = 0; #10;
    a = 1; b = 0; c = 0; d = 1; #10;
    a = 1; b = 0; c = 1; d = 0; #10;
    a = 1; b = 0; c = 1; d = 1; #10;
    a = 1; b = 1; c = 0; d = 0; #10;
    a = 1; b = 1; c = 0; d = 1; #10;
    a = 1; b = 1; c = 1; d = 0; #10;
    a = 1; b = 1; c = 1; d = 1; #10;


    $display("complete!!!");

end

endmodule
